`timescale 1ns / 1ps



module Syndrome(    
        input  R,
        input CLK,          
        input reset,
        output reg [16199:0] Cfront=0,
        //output enerror,            �Ȳ�Ҫ��  2019.05.26
        
        output reg enableBM=0,//    2019/5/25 �¼ӵ�
        
                   output reg [15:0] S1=0,    //У���ӼĴ���
                   output reg [15:0] S2=0,
                   output reg [15:0] S3=0,
                   output reg [15:0] S4=0,
                   output reg[15:0] S5=0,
                   output reg[15:0] S6=0,
                   output reg[15:0] S7=0,
                   output reg[15:0] S8=0,
                   output reg[15:0] S9=0,
                   output reg[15:0] S10=0,
                   output reg[15:0] S11=0,
                   output reg[15:0] S12=0,
                   output reg[15:0] S13=0,     
                   output reg[15:0] S14=0,
                   output reg[15:0] S15=0,
                   output reg[15:0] S16=0,
                   output reg[15:0] S17=0,
                   output reg[15:0] S18=0,
                   output reg[15:0] S19=0,
                   output reg[15:0] S20=0,
                   output reg[15:0] S21=0,
                   output reg[15:0] S22=0,
                   output reg[15:0] S23=0
        
        );
           
           //reg [195:0]controlg=196'ha7130741c22e288e2867966c6e1a844481a3c2fbb3012af38;
           reg [16:0]g1=17'd65581;      
           reg [16:0]g2=17'd65907;
           reg [16:0]g3=17'd69565;
           reg [16:0]g4=17'd88629;
           reg [16:0]g5=17'd73503;
           reg [16:0]g6=17'd128949;
           reg [16:0]g7=17'd110437;
           reg [16:0]g8=17'd95079;
           reg [16:0]g9=17'd95655;
           reg [16:0]g10=17'd80429;
           reg [16:0]g11=17'd65907;
           reg [16:0]g12=17'd72419;
           
          
           
           reg [15:0]b1=0;               //12��������·�ֱ�ļĴ��������Ǽ���У���ӵ�ri
           reg [15:0]b2=0;
           reg [15:0]b3=0;
           reg [15:0]b4=0;
           reg [15:0]b5=0;
           reg [15:0]b6=0;
           reg [15:0]b7=0;
           reg [15:0]b8=0;
           reg [15:0]b9=0;
           reg [15:0]b10=0;
           reg [15:0]b11=0;
           reg [15:0]b12=0;
           
           reg [11:0]b16=0;      //linshicunfangzuigaowei   ��ʱ������λ
           reg [3:0]ib16=0;      //b16 de xunhuanbianliang,bazhishuchugei12gechufadianlu   
           
           
           
                  
           //reg [191:0]Bbs=0;                                 //    ���ڽ���֮�����µľ���ϵ��ri
           //reg inputdata=0;
           reg [14:0]count=0;
           reg [4:0]i=0;                 //yonglaigeimeige chufadianlude jicunqi fuzhide
           reg b191=0;
           reg [7:0] j=191;
           reg midd;
           

           
           
           always@(posedge CLK  or negedge reset)    
              begin
              if (!reset)//if(!a)�������aΪ�棬Ҳ����aΪ0ʱ��if������������֮��������
              begin
              //Bbs=0;
              
              
              b1=0;
              b2=0;
              b3=0;
              b4=0;
              b5=0;
              b6=0;
              b7=0;
              b8=0;
              b9=0;
              b10=0;
              b11=0;
              b12=0;
              
              ib16=0;
              
              end
              count=count+1;
              //bits=Bbs;
              
              if (count<=16200)                                         //16200������������
                 begin
                    //inputdata<={$random} % 2;
                    //dataout=R;                                 xianbushuchu
                    
                    if (count<=16008)
                    Cfront[count-1]=R;                                //ֱ�Ӵ�Ž��յ�����   2019.05.26��һ��always
                    
                    for (ib16=0; ib16<=11 ; ib16=ib16+1)            //12��������·��
                    begin
                    case(ib16)
                    0:begin                    b16[0]=b1[15];                                  b1=b1<<1;             b1[0]=R^b1[15];
                                           for( i=1 ; i<=15 ; i=i+1 )                //
                                           begin
                                                                   
                                           b1[i]=b1[i]^(g1[i]&b1[0]);   //haoxiangmeiyunxing
                                              
                                           end    
                    
                    
                                         end
                    1:begin                    b16[1]=b2[15];                                  b2=b2<<1;               b2[0]=R^b2[15];    
                                                          for( i=1 ; i<=15 ; i=i+1 )                //
                                                          begin
                                                                                  
                                                          b2[i]=b1[i]^(g2[i]&b2[0]);   //haoxiangmeiyunxing
                                                             
                                                          end    
                                     end   
                    2:begin                    b16[2]=b3[15];                                  b3=b3<<1;               b3[0]=R^b3[15];   
                                                          for( i=1 ; i<=15 ; i=i+1 )                //
                                                          begin
                                                                                  
                                                          b3[i]=b3[i]^(g3[i]&b3[0]);   //haoxiangmeiyunxing
                                                             
                                                          end    
                                                                           end
                    3:begin                    b16[3]=b4[15];                                  b4=b4<<1;               b4[0]=R^b4[15];           
                                                          for( i=1 ; i<=15 ; i=i+1 )                //
                                                          begin
                                                                                  
                                                          b4[i]=b4[i]^(g4[i]&b4[0]);   //haoxiangmeiyunxing
                                                             
                                                          end    
                            end
                    4:begin                    b16[4]=b5[15];                                  b5=b5<<1;               b5[0]=R^b5[15];        
                                                          for( i=1 ; i<=15 ; i=i+1 )                //
                                                          begin
                                                                                  
                                                          b5[i]=b5[i]^(g5[i]&b5[0]);   //haoxiangmeiyunxing
                                                             
                                                          end    
                                                                    end
                    5:begin                    b16[5]=b6[15];                                  b6=b6<<1;               b6[0]=R^b6[15];        
                                                          for( i=1 ; i<=15 ; i=i+1 )                //
                                                          begin
                                                                                  
                                                          b6[i]=b6[i]^(g6[i]&b6[0]);   //haoxiangmeiyunxing
                                                             
                                                          end    
                              end
                    6:begin                    b16[6]=b7[15];                                  b7=b7<<1;               b7[0]=R^b7[15];           
                                                          for( i=1 ; i<=15 ; i=i+1 )                //
                                                          begin
                                                                                  
                                                          b7[i]=b7[i]^(g7[i]&b7[0]);   //haoxiangmeiyunxing
                                                             
                                                          end    
                           end
                    7:begin                    b16[7]=b8[15];                                  b8=b8<<1;               b8[0]=R^b8[15];        
                                                          for( i=1 ; i<=15 ; i=i+1 )                //
                                                          begin
                                                                                  
                                                          b8[i]=b8[i]^(g8[i]&b8[0]);   //haoxiangmeiyunxing
                                                             
                                                          end    
                              end
                    8:begin                    b16[8]=b9[15];                                  b9=b9<<1;               b9[0]=R^b9[15];           
                                                          for( i=1 ; i<=15 ; i=i+1 )                //
                                                          begin
                                                                                  
                                                          b9[i]=b9[i]^(g9[i]&b9[0]);   //haoxiangmeiyunxing
                                                             
                                                          end    
                             end
                    9:begin                    b16[9]=b10[15];                                 b10=b10<<1;             b10[0]=R^b10[15];         
                     for( i=1 ; i<=15 ; i=i+1 )                //
                                                          begin
                                                                                  
                                                          b10[i]=b10[i]^(g10[i]&b10[0]);   //haoxiangmeiyunxing
                                                             
                                                          end    
                                                                      end
                    10:begin                   b16[10]=b11[15];                                b11=b11<<1;            b11[0]=R^b11[15];       
                                                          for( i=1 ; i<=15 ; i=i+1 )                //
                                                          begin
                                                                                  
                                                          b11[i]=b11[i]^(g11[i]&b11[0]);   //haoxiangmeiyunxing
                                                             
                                                          end    
                                 end
                    11:begin                   b16[11]=b12[15];                                b12=b12<<1;            b12[0]=R^b12[15];      
                                                          for( i=1 ; i<=15 ; i=i+1 )                //
                                                          begin
                                                                                  
                                                          b12[i]=b12[i]^(g12[i]&b12[0]);   //haoxiangmeiyunxing
                                                             
                                                          end    
                                 end
                                   
                    
                    endcase
                  end
                    
                    
              end              //line 80   'if'               //shurudexiancunqilai
                    /*         b191=Bbs[191];                        //liuyiweicunfangyiweidegaowei
                    Bbs=Bbs<<1;        //
                    Bbs[0]=b191^R;                   
                     for( i=1 ; i<=191 ; i=i+1 )                //
                            begin
                                                    
                            Bbs[i]=Bbs[i]^(controlg[i+3]&Bbs[0]);   //haoxiangmeiyunxing
                               
                            end    
       //��ѭ��
                 end                          */
        /*      else if (count<=16200&&count>=16009)
                  begin 
                     dataout=Bbs[j];
                     j=j-1;  
                  end                 */
            if (count==16200)     
                  begin                  //֮���synchronized �����ȫ���ƹ���
          S1[15]=b1[15]; 
                  S1[14]=b1[14];
                  S1[13]=b1[13];
                  S1[12]=b1[12];
                  S1[11]=b1[11];
                  S1[10]=b1[10];
                  S1[9]=b1[9];
                  S1[8]=b1[8];
                  S1[7]=b1[7];
                  S1[6]=b1[6];
                  S1[5]=b1[5];
                  S1[4]=b1[4];
                  S1[3]=b1[3];
                  S1[2]=b1[2];
                  S1[1]=b1[1];
                  S1[0]=b1[0];
                  
                  S2[15]=b1[13]^b1[14];
                  S2[14]=b1[15]^b1[14]^b1[7];
                  S2[13]=b1[12] ^ b1[13];
                  S2[12]=b1[6] ^ b1[13] ^ b1[14];
                  S2[11]=b1[11] ^ b1[12];
                  S2[10]=b1[5] ^b1[12] ^ b1[13];
                  S2[9]=b1[10] ^ b1[11];
                  S2[8]=b1[4]^ b1[11] ^ b1[12] ^ b1[15];
                  S2[7]=b1[9] ^ b1[10];
                  S2[6]=b1[3] ^ b1[10] ^ b1[11] ^ b1[14];
                  S2[5]=b1[8] ^ b1[9];
                  S2[4]=b1[2] ^ b1[9] ^ b1[10] ^ b1[14] + b1[15];
                  S2[3]=b1[8] ^ b1[14] ^ b1[15];
                  S2[2]=b1[1] ^ b1[8] ^ b1[9] ^ b1[15];
                  S2[1]=b1[14] ^ b1[15]; 
                  S2[0]=b1[0] ^ b1[8] ^ b1[15];
                  
                  
                  S3[15]=b2[5];
                  S3[14]=b2[12]^b2[14]^b2[10]^b2[9];// r9 + r10 + r12 + r14
                  S3[13]=b2[15]^b2[13]^b2[9]^b2[8];// r8 + r9 + r13 + r15,
                  S3[12]=b2[15]^b2[4];// r4 + r15,
                  S3[11]=b2[13]^b2[11]^b2[9]^b2[8];//r8 + r9 + r11 + r13,
                  S3[10]=b2[15]^b2[14]^b2[12]^b2[8]^b2[7];//r7 + r8 + r12 + r14 + r15,
                  S3[9]=b2[15]^b2[14]^b2[3];//r3 + r14 + r15,
                  S3[8]=b2[15]^b2[12]^b2[10]^b2[8]^b2[7];//r7 + r8 + r10 + r12 + r15,
                  S3[7]=b2[15]^b2[14]^b2[13]^b2[11]^b2[6]^b2[7];//r6 + r7 + r11 + r13 + r14 + r15,
                  S3[6]=b2[13]^b2[14]^b2[2];//r2 + r13 + r14,
                  S3[5]=b2[15]^b2[14]^b2[11]^b2[7]^b2[9]^b2[6];//r6 + r7 + r9 + r11 + r14 + r15,
                  S3[4]=b2[13]^b2[14]^b2[15]^b2[12]^b2[10]^b2[6];//r6 + r10 + r12 + r13 + r14 + r15,
                  S3[3]=b2[13]^b2[14]^b2[10]^b2[9]^b2[1];                     // r1 + r9 + r10 + r13 + r14,
                  S3[2]=b2[10]^b2[14]^b2[6]^b2[9];//r6 + r9 + r10 + r14,
                  S3[1]=b2[13]^b2[15]^b2[10]^b2[11];                                //r10 + r11 + r13 + r15,
                  S3[0]=b2[14]^b2[10]^b2[0]^b2[9];//r0 + r9 + r10 + r14,
                  
                  
                                S4[15]=b1[15]^b1[14]^b1[12] ^ b1[13]^b1[7];//r7 + r12 + r13 + r14 + r15,
                                S4[14]=b1[15]^b1[13]^b1[10]^b1[9]^b1[7];//r7 + r9 + r10 + r13 + r15, 
                                S4[13]=b1[12] ^ b1[14]^b1[6];// r6 + r12 + r14,
                                S4[12]=b1[15]^b1[13]^b1[12]^b1[11]^b1[10]^b1[3]^b1[7];//r3 + r7 + r10 + r11 + r12 + r13 + r15, 
                                S4[11]=b1[11] ^ b1[14]^b1[12] ^ b1[13]^b1[6];//r6 + r11 + r12 + r13 + r14,
                                S4[10]=b1[6]^b1[8]^b1[9] ^b1[12] ^ b1[14];//r6 + r8 + r9 + r12 + r14,
                                S4[9]=b1[5]^b1[11] ^ b1[13];//r5 + r11 + r13,
                                S4[8]=b1[2]^b1[6]^b1[9]^b1[10]^ b1[11] ^ b1[12] ^b1[14]^ b1[15];//r2 + r6 + r9 + r10 + r11 + r12 + r14 + r15,
                                S4[7]=b1[5]^b1[11] ^ b1[13]^b1[12] ^ b1[10];//r5 + r10 + r11 + r12 + r13,
                                S4[6]=b1[5]^b1[7]^b1[8]^b1[11] ^ b1[13];//r5 + r7 + r8 + r11 + r13,
                                S4[5]=b1[4] ^b1[10]^b1[12] ^ b1[15];//r4 + r10 + r12 + r15,
                                S4[4]=b1[1]^b1[5] ^ b1[7] ^ b1[8] ^ b1[9] ^ b1[10] ^b1[11] ^ b1[12];// r1 + r5 + r7 + r8 + r9 + r10 + r11 + r12,
                                S4[3]=b1[7] ^ b1[4] ^b1[11]^b1[12] ^ b1[13];//r4 + r7 + r11 + r12 + r13,
                                S4[2]=b1[4] ^ b1[10] ^ b1[12] ^ b1[13];//r4 + r10 + r12 + r13,
                                S4[1]=b1[13] ^ b1[15]^b1[7]; //r7 + r13 + r15, 
                                S4[0]=b1[0] ^ b1[8] ^b1[4] ^b1[11]^b1[12] ^ b1[13]^ b1[14];//r0 + r4 + r8 + r11 + r12 + r13 + r14,
                
                
                
                
                                                           S5[15]=b3[15]^b3[14]^b3[12]^b3[11]^b3[10]^b3[3];// r3 + r10 + r11 + r12 + r14 + r15,
                                                           S5[14]=b3[5]^b3[6]^b3[14]^b3[12]^b3[11]^b3[10]^b3[8];// r5 + r6 + r8 + r10 + r11 + r12 + r14,
                                                           S5[13]=b3[13]^b3[14]^b3[7]^b3[10]^b3[9];//  r7 + r9 + r10 + r13 + r14,
                                                           S5[12]=b3[15]^b3[9]^b3[14]^b3[12]^b3[11]^b3[10]^b3[8]^b3[5];// r5 + r8 + r9 + r10 + r11 + r12 + r14 + r15,
                                                           S5[11]=b3[15]^b3[5];//r5 + r15,
                                                           S5[10]=b3[2]^b3[15]^b3[14]^b3[13]^b3[11]^b3[10]^b3[9];//r2 + r9 + r10 + r11 + r13 + r14 + r15,
                                                           S5[9]=b3[4]^b3[5]^b3[7]^b3[9]^b3[10]^b3[11]^b3[13];//r4 + r5 + r7 + r9 + r10 + r11 + r13,
                                                           S5[8]=b3[15]^b3[13]^b3[12]^b3[9]^b3[8]^b3[6];//r6 + r8 + r9 + r12 + r13 + r15,
                                                           S5[7]=b3[15]^b3[14]^b3[13]^b3[11]^b3[10]^b3[9]^b3[8]^b3[7]^b3[4];//r4 + r7 + r8 + r9 + r10 + r11 + r13 + r14 + r15,
                                                           S5[6]=b3[4]^b3[14]^b3[15];//r4 + r14 + r15,
                                                           S5[5]=b3[1] ^b3[8]^b3[9]^b3[14]^b3[12]^b3[13]^b3[10];// r1 + r8 + r9 + r10 + r12 + r13 + r14,
                                                           S5[4]=b3[4]^b3[15]^b3[14]^b3[9]^b3[11]^b3[8]^b3[6];//   r4 + r6 + r8 + r9 + r11 + r14 + r15,
                                                           S5[3]=b3[7] ^b3[6]^b3[10];//  r6 + r7 + r10,
                                                           S5[2]=b3[15]^b3[14]^b3[8]^b3[11]^b3[10]^b3[6];//    r6 + r8 + r10 + r11 + r14 + r15,
                                                           S5[1]=b3[13]^b3[15]^b3[9]^b3[12]^b3[11]^b3[10]^b3[6]; //   r6 + r9 + r10 + r11 + r12 + r13 + r15,
                                                           S5[0]=b3[0]^ b3[6];//            r0 + r6,
                  
                  
                  
                  
                                                                        S6[15]=b2[15]^b2[14]^b2[13]^b2[12]^b2[10]^b2[8];//     r8 + r10 + r12 + r13 + r14 + r15,
                                                                        S6[14]=b2[15]^b2[13]^b2[12]^b2[11]^b2[10]^b2[9]^b2[6]^b2[7]^b2[5];//    r5 + r6 + r7 + r9 + r10 + r11 + r12 + r13 + r15, 
                                                                        S6[13]=b2[4]^b2[13]^b2[9]^b2[8];//         r4 + r8 + r9 + r13,
                                                                        S6[12]=b2[15]^b2[2]^b2[12]^b2[10]^b2[8];//              r2 + r8 + r10 + r12 + r15,
                                                                        S6[11]=b2[15]^b2[4]^b2[9]^b2[11]^b2[13]^b2[8];//            r4 + r8 + r9 + r11 + r13 + r15,
                                                                        S6[10]=b2[6]^b2[4]^b2[15]^b2[14]^b2[13]^b2[11]^b2[8]^b2[7];// r4 + r6 + r7 + r8 + r11 + r13 + r14 + r15,
                                                                        S6[9]=b2[15]^b2[14]^b2[7]^b2[11]^b2[13]^b2[12]^b2[9];//         r7 + r9 + r11 + r12 + r13 + r14 + r15,
                                                                        S6[8]=b2[14]^b2[12]^b2[11]^b2[10]^b2[9]^b2[6]^b2[5]^b2[4]^b2[8];//r4 + r5 + r6 + r8 + r9 + r10 + r11 + r12 + r14,
                                                                        S6[7]=b2[3]^b2[8]^b2[12]^b2[7];//                r3 + r7 + r8 + r12,
                                                                        S6[6]=b2[15]^b2[14]^b2[11]^b2[9]^b2[7]^b2[1];//          r1 + r7 + r9 + r11 + r14 + r15,
                                                                        S6[5]=b2[14]^b2[12]^b2[10]^b2[8]^b2[7]^b2[3];//           r3 + r7 + r8 + r10 + r12 + r14,
                                                                        S6[4]=b2[8]^b2[7]^b2[6]^b2[5]^b2[3];//                      r3 + r5 + r6 + r7 + r8,
                                                                        S6[3]=b2[15]^b2[14]^b2[9]^b2[8]^b2[7]^b2[5];                     //                r5 + r7 + r8 + r9 + r14 + r15,  
                                                                        S6[2]=b2[15]^b2[14]^b2[13]^b2[12]^b2[11]^b2[8]^b2[7]^b2[5]^b2[3];//r3 + r5 + r7 + r8 + r11 + r12 + r13 + r14 + r15,
                                                                        S6[1]=b2[14]^b2[12]^b2[10]^b2[9]^b2[5];                                //               r5 + r9 + r10 + r12 + r14,
                                                                        S6[0]=b2[15]^b2[14]^b2[12]^b2[9]^b2[8]^b2[7]^b2[5]^b2[0];//          r0 + r5 + r7 + r8 + r9 + r12 + r14 + r15,
                  
                  
                                                               S7[15]=b4[15]^b4[13]^b4[12]^b4[11]^b4[10]^b4[9]^b4[8]^b4[4];//     r4 + r8 + r9 + r10 + r12 + r13 + r15,
                                                               S7[14]=b4[15]^b4[14]^b4[11]^b4[10]^b4[7]^b4[6]^b4[4]^b4[2];//     r2 + r4 + r6 + r7 + r10 + r11 + r14 + r15,
                                                               S7[13]=b4[13]^b4[11]^b4[10]^b4[8]^b4[7]^b4[5];//                  r5 + r7 + r8 + r10 + r11 + r13,
                                                               S7[12]=b4[14]^b4[13]^b4[11]^b4[10]^b4[7]^b4[8]^b4[5];//                   r4 + r7 + r10 + r11 + r13 + r14,
                                                               S7[11]=b4[15]^b4[13]^b4[9]^b4[8]^b4[7];//               r7 + r8 + r9 + r13 + r15,
                                                               S7[10]=b4[15]^b4[13]^b4[12]^b4[11]^b4[10]^b4[6]^b4[8]^b4[3];//         r3 + r6 + r8 + r10 + r11 + r12 + r13 + r15,
                                                               S7[9]=b4[15]^b4[14]^b4[12]^b4[11]^b4[7]^b4[6]^b4[5];//         r5 + r6 + r7 + r11 + r12 + r14 + r15, 
                                                               S7[8]=b4[15]^b4[14]^b4[12]^b4[11]^b4[7]^b4[9]^b4[8]^b4[3];//        r3 + r7 + r8 + r9 + r11 + r12 + r14 + r15,
                                                               S7[7]=b4[15]^b4[13]^b4[14]^b4[6]^b4[10]^b4[9]^b4[5]^b4[3]^b4[1];//               r1 + r3 + r5 + r6 + r9 + r10 + r13 + r14 + r15,
                                                               S7[6]=b4[15]^b4[12]^b4[4]^b4[10]^b4[9]^b4[7]^b4[6];//           r4 + r6 + r7 + r9 + r10 + r12 + r15,
                                                               S7[5]=b4[15]^b4[13]^b4[12]^b4[10]^b4[9]^b4[6]^b4[3];//            r3 + r6 + r9 + r10 + r12 + r13 + r15,
                                                               S7[4]=b4[14]^b4[13]^b4[10]^b4[9]^b4[7]^b4[6]^b4[4];//                      r4 + r6 + r7 + r9 + r10 + r13 + r14,
                                                               S7[3]=b4[12]^b4[10]^b4[9]^b4[6]^b4[5]^b4[4];                     //                    r4 + r5 + r6 + r9 + r12,       
                                                               S7[2]=b4[15]^b4[14]^b4[13]^b4[12]^b4[10]^b4[9]^b4[7]^b4[6];//       r6 + r7 + r9 + r10 + r12 + r13 + r14 + r15,
                                                               S7[1]=b4[14]^b4[13]^b4[12]^b4[11]^b4[9]^b4[7]^b4[6];              //                r4 + r7 + r9 + r11 + r12 + r13 + r14,
                                                               S7[0]=b4[15]^b4[13]^b4[12]^b4[8]^b4[7]^b4[6]^b4[0];//              r0 + r6 + r7 + r8 + r12 + r13 + r15,
                  
                  
        
         S8[15]=b1[15]^b1[14]^b1[13]^b1[12]^b1[7];//r6 + r7 + r9 + r10 + r12 + r13 + r14 + r15,
         S8[14]=b1[15]^b1[13]^b1[10]^b1[9]^b1[7];//               r5 + r9 + r11 + r13 + r14,
         S8[13]=b1[12] ^ b1[14]^b1[6];//     r3 + r6 + r7 + r10 + r11 + r13 + r14 + r15,
         S8[12]=b1[15]^b1[13]^b1[12]^b1[11]^b1[10]^b1[3]^b1[7];//   r5 + r6 + r8 + r9 + r10 + r11 + r12 + r14 + r15,
         S8[11]=b1[11] ^ b1[14]^b1[12] ^ b1[13]^b1[6];//         r3 + r6 + r7 + r10 + r14 + r15,
         S8[10]=b1[6]^b1[8]^b1[9] ^b1[12] ^ b1[14];//     r3 + r4 + r6 + r7 + r11 + r12 + r13 + r14,
         S8[9]=b1[5]^b1[11] ^ b1[13];//                          r8 + r9 + r11 + r13,
         S8[8]=b1[2]^b1[6]^b1[9]^b1[10]^ b1[11] ^ b1[12] ^b1[14]^ b1[15];//    r1 + r3 + r5 + r6 + r7 + r8 + r9 + r11 + r13
         S8[7]=b1[5]^b1[11] ^ b1[13]^b1[12] ^ b1[10];//      r5 + r6 + r8 + r9 + r11 + r12 + r13 + r14,
         S8[6]=b1[5]^b1[7]^b1[8]^b1[11] ^ b1[13];//  r4 + r8 + r10 + r12 + r13 + r15,
         S8[5]=b1[4] ^b1[10]^b1[12] ^ b1[15];//  r2 + r5 + r6 + r9 + r10 + r12 + r13 + r14 + r15,
         S8[4]=b1[1]^b1[5] ^ b1[7] ^ b1[8] ^ b1[9] ^ b1[10] ^b1[11] ^ b1[12];//            r4 + r5 + r6 + r8 + r11 + r12,
         S8[3]=b1[7] ^ b1[4] ^b1[11]^b1[12] ^ b1[13];// r2 + r6 + r11 + r15,
         S8[2]=b1[4] ^ b1[10] ^ b1[12] ^ b1[13];//  r2 + r5 + r6 + r9 + r10 + r13 + r15,
         S8[1]=b1[13] ^ b1[15]^b1[7]; //               r9 + r10 + r12 + r14,
         S8[0]=b1[0] ^ b1[8] ^b1[4] ^b1[11]^b1[12] ^ b1[13]^ b1[14];// r0 + r2 + r4 + r6 + r7 + r8 + r9 + r10 + r12 + r14,
        
        
        
         S9[15]=b5[7]^b5[8]^b5[10]^b5[11]^b5[13];                         //r7 + r8 + r10 + r11 + r13,
         S9[14]=b5[3]^b5[4]^b5[6]^b5[8]^b5[9]^b5[10]^b5[12]^b5[15];//              r3 + r4 + r6 + r8 + r9 + r10 + r12 + r15,
         S9[13]=b5[3]^b5[5]^b5[6]^b5[9]^b5[11]^b5[12];//      r3 + r5 + r6 + r9 + r11 + r12,
         S9[12]=b5[5]^b5[8]^b5[9]^b5[10]^b5[12]^b5[13]^b5[14];//       r5 + r8 + r9 + r10 + r12 + r13 + r14,
         S9[11]=b5[3]^b5[6]^b5[7]^b5[10]^b5[12]^b5[14]^b5[15];//               r3 + r6 + r7 + r10 + r12 + r14 + r15,
         S9[10]=b5[4]^b5[5]^b5[10]^b5[11]^b5[12]^b5[13]^b5[14];//              r4 + r5 + r10 + r11 + r12 + r13 + r14, 
         S9[9]=b5[1]^b5[5]^b5[6]^b5[8]^b5[10]^b5[11]^b5[12]^b5[13]^b5[14]^b5[15];//                         r1 + r5 + r6 + r8 + r10 + r11 + r12 + r13 + r14 + r15, 
         S9[8]=b5[4]^b5[5]^b5[6]^b5[7]^b5[8]^b5[11]^b5[12]^b5[13]^b5[14];//          r4 + r5 + r6 + r7 + r8 + r11 + r12 + r13 + r14,
         S9[7]=b5[2]^b5[5]^b5[7]^b5[8]^b5[9]^b5[12]^b5[15];//                  r2 + r5 + r7 + r8 + r9 + r12 + r15,  
         S9[6]=b5[6]^b5[7]^b5[9]^b5[10]^b5[12]^b5[15];//                  r6 + r7 + r9 + r10 + r12 + r15,
         S9[5]=b5[2]^b5[3]^b5[5]^b5[7]^b5[8]^b5[9]^b5[11]^b5[14]^b5[15];//         r2 + r3 + r5 + r7 + r8 + r9 + r11 + r14 + r15,
         S9[4]=b5[2]^b5[4]^b5[7]^b5[13]^b5[15];//                   r2 + r4 + r5 + r7 + r13 + r15,
         S9[3]=b5[3]^b5[4]^b5[6]^b5[7]^b5[10]^b5[11]^b5[13];//               r3 + r6 + r7 + r10 + r11 + r13,
         S9[2]=b5[2]^b5[3]^b5[7]^b5[8]^b5[10]^b5[11]^b5[12]^b5[14]^b5[15];//     r2 + r3 + r7 + r8 + r10 + r11 + r12 + r14 + r15,
         S9[1]=b5[5]^b5[6]^b5[7]^b5[8]^b5[9]^b5[12]^b5[13]^b5[14]^b5[15]; //                 r5 + r6 + r7 + r8 + r9 + r12 + r13 + r14 + r15,
         S9[0]=b5[0]^b5[3]^b5[6]^b5[8]^b5[9]^b5[10]^b5[13];//           r0 + r3 + r6 + r8 + r9 + r10 + r13,              
                  
         S10[15]=b3[5]^b3[6]^b3[7]^b3[8]^b3[9]^b3[11]^b3[12]^b3[13];//                 r5 + r6 + r7 + r8 + r9 + r11 + r12 + r13,
         S10[14]=b3[3]^b3[4]^b3[5]^b3[6]^b3[7]^b3[9]^b3[10]^b3[11]^b3[13]^b3[14];//            r3 + r4 + r5 + r6 + r7 + r9 + r10 + r11 + r13 + r14,
         S10[13]=b3[5]^b3[7]^b3[8]^b3[11]^b3[12]^b3[13]^b3[15];//    r5 + r7 + r8 + r11 + r12 + r13 + r15,
         S10[12]=b3[4]^b3[5]^b3[6]^b3[7]^b3[8]^b3[9]^b3[11]^b3[12]^b3[13]^b3[14]^b3[15];//       r4 + r5 + r6 + r7 + r8 + r9 + r11 + r12 + r13 + r14 + r15,
         S10[11]=b3[8]^b3[9]^b3[10]^b3[11]^b3[12]^b3[14];                    //               r8 + r9 + r10 + r11 + r12 + r14,
         S10[10]=b3[1]^b3[5]^b3[7]^b3[9]^b3[10]^b3[11]^b3[14]^b3[15];//            r1 + r5 + r7 + r9 + r10 + r11 + r14 + r15,
         S10[9]=b3[2]^b3[5]^b3[9]^b3[10]^b3[11]^b3[13]^b3[14];//                 r2 + r5 + r9 + r10 + r11 + r13 + r14,
         S10[8]=b3[3]^b3[4]^b3[6]^b3[11]^b3[14];//                             r3 + r4 + r6 + r11 + r14,
         S10[7]=b3[2]^b3[4]^b3[5]^b3[7]^b3[14]^b3[15];//           r2 + r4 + r5 + r7 + r14 + r15,
         S10[6]=b3[2]^b3[7]^b3[8]^b5[9]^b3[10]^b3[12]^b3[13];//                r2 + r7 + r8 + r9 + r10 + r12 + r13,
         S10[5]=b3[4]^b3[5]^b3[6]^b3[7]^b3[8]^b3[10]^b3[11]^b3[12]^b3[15];//              r4 + r5 + r6 + r7 + r8 + r10 + r11 + r12 + r15,
         S10[4]=b3[2]^b3[3]^b3[4]^b3[7]^b3[10]^b3[11]^b3[15];//                           r2 + r3 + r4 + r7 + r10 + r11 + r15,
         S10[3]=b3[3]^b3[5]^b3[9]^b3[12]^b3[13];//                  r3 + r5 + r9 + r12 + r13,
         S10[2]=b3[3]^b3[4]^b3[5]^b3[7]^b3[8]^b3[9]^b3[10]^b3[11]^b3[12]^b3[13]^b3[14]^b3[15];//    r3 + r4 + r5 + r7 + r8 + r9 + r10 + r11 + r12 + r13 + r14 + r15,
         S10[1]=b3[3]^b3[5]^b3[6]^b3[8]^b3[15]; //                  r3 + r5 + r6 + r8 + r15, 
         S10[0]=b3[0]^b3[3]^b3[8]^b3[9]^b3[10]^b3[11]^b3[13]^b3[14];//                        r0 + r3 + r8 + r9 + r10 + r11 + r13 + r14,  
         
         
         S11[15]=b6[5]^b6[9]^b6[10]^b6[12]^b6[13]^b6[15];//                 r5 + r9 + r10 + r12 + r13 + r15,
         S11[14]=b6[5]^b6[6]^b6[7]^b6[8]^b6[10]^b6[11]^b6[12]^b6[13]^b6[14]^b6[15];//          r5 + r6 + r7 + r8 + r10 + r11 + r12 + r13 + r14 + r15,
         S11[13]=b6[7]^b6[8]^b6[9]^b6[10]^b6[11]^b6[13]^b6[15];//              r7 + r8 + r9 + r10 + r11 + r13 + r15,
         S11[12]=b6[4]^b6[5]^b6[7]^b6[8]^b6[10]^b6[11]^b6[13];//               r4 + r5 + r7 + r8 + r10 + r11 + r13,
         S11[11]=b6[1]^b6[2]^b6[3]^b6[4]^b6[6]^b6[10]^b6[12]^b6[13]^b6[14]^b6[15];           //            r1 + r2 + r3 + r4 + r6 + r10 + r12 + r13 + r14 + r15,
         S11[10]=b6[5]^b6[6]^b6[7]^b6[8]^b6[9]^b6[10]^b6[13];//                r5 + r6 + r7 + r8 + r9 + r10 + r13,
         S11[9]=b6[2]^b6[4]^b6[5]^b6[6]^b6[7]^b6[8]^b6[9]^b6[10]^b6[14]^b6[15];//                r2 + r4 + r5 + r6 + r7 + r8 + r9 + r10 + r14 + r15,,
         S11[8]=b6[2]^b6[4]^b6[6]^b6[7]^b6[8]^b6[9]^b6[10]^b6[12]^b6[14];//                         r2 + r4 + r6 + r7 + r8 + r9 + r10 + r12 + r14,
         S11[7]=b6[3]^b6[4]^b6[5]^b6[8]^b6[11]^b6[15];//                  r3 + r4 + r5 + r8 + r11 + r15,
         S11[6]=b6[2]^b6[4]^b6[6]^b6[11]^b6[12]^b6[13]^b6[15];//                   r2 + r4 + r6 + r11 + r12 + r13 + r15,
         S11[5]=b6[3]^b6[9]^b6[10]^b6[11]^b6[13]^b6[14]^b6[15];//                 r3 + r9 + r10 + r11 + r13 + r15, 
         S11[4]=b6[4]^b6[5]^b6[8]^b6[10]^b6[11]^b6[13]^b6[14]^b6[15];//                        r4 + r5 + r8 + r10 + r11 + r13 + r14 + r15,
         S11[3]=b6[4]^b6[8]^b6[9]^b6[15];//                         r4 + r8 + r9 + r15,
         S11[2]=b6[5]^b6[6]^b6[9]^b6[10]^b6[11]^b6[14];//    r5 + r6 + r9 + r10 + r11 + r14,
         S11[1]=b6[3]^b6[5]^b6[7]^b6[12]^b6[13]^b6[14]; //                   r3 + r5 + r7 + r12 + r13 + r14,
         S11[0]=b6[0]^b6[4]^b6[10]^b6[11]^b6[12]^b6[14];//                             r0 + r4 + r10 + r11 + r12 + r14,           
         
         
         S12[15]=b2[4]^b2[5]^b2[6]^b2[7]^b2[8]^b2[10]^b2[11]^b2[12]^b2[15];           //   r4 + r5 + r6 + r7 + r8 + r10 + r11 + r12 + r15,
         S12[14]=b2[3]^b2[5]^b2[6]^b2[9]^b2[11]^b2[12]^b2[14];//       r3 + r5 + r6 + r9 + r11 + r12 + r14,
         S12[13]=b2[2]^b2[4]^b2[9]^b2[10]^b2[12]^b2[13]^b2[15];//          r2 + r4 + r9 + r10 + r12 + r13 + r15,
         S12[12]=b2[1]^b2[4]^b2[5]^b2[6]^b2[8]^b2[9]^b2[10]^b2[12]^b2[14];//               r1 + r4 + r5 + r6 + r8 + r9 + r10 + r12 + r14,
         S12[11]=b2[2]^b2[4]^b2[9]^b2[10]^b2[11]^b2[12]^b2[13];//      r2 + r4 + r9 + r10 + r11 + r12 + r13,
         S12[10]=b2[2]^b2[3]^b2[4]^b2[7]^b2[8]^b2[9]^b2[13]^b2[14]^b2[15];//    r2 + r3 + r4 + r7 + r8 + r9 + r13 + r14 + r15,
         S12[9]=b2[6]^b2[7]^b2[9]^b2[14];//         r6 + r7 + r9 + r14,
         S12[8]=b2[2]^b2[3]^b2[4]^b2[5]^b2[6]^b2[7]^b2[9]^b2[11]^b2[14]^b2[15];// r2 + r3 + r4 + r5 + r6 + r7 + r9 + r11 + r14 + r15,
         S12[7]=b2[4]^b2[6]^b2[8]^b2[9]^b2[12];//       r4 + r6 + r8 + r9 + r12,
         S12[6]=b2[7]^b2[8]^b2[9]^b2[10]^b2[11]^b2[12]^b2[13];//            r7 + r8 + r9 + r10 + r11 + r12 + r13,
         S12[5]=b2[4]^b2[5]^b2[6]^b2[7]^b2[8]^b2[10]^b2[13]^b2[15];//       r4 + r5 + r6 + r7 + r8 + r10 + r13 + r15,
         S12[4]=b2[3]^b2[4]^b2[8]^b2[13]^b2[15];//         r3 + r4 + r8 + r13 + r15,
         S12[3]=b2[4]^b2[7]^b2[10]^b2[12];                     //             r4 + r7 + r10 + r12,
         S12[2]=b2[4]^b2[6]^b2[7]^b2[9]^b2[10];//               r4 + r6 + r7 + r9 + r10,
         S12[1]=b2[5]^b2[6]^b2[7]^b2[8]^b2[9]^b2[11]^b2[14];                                //     r5 + r6 + r7 + r8 + r9 + r11 + r14,
         S12[0]=b2[0]^b2[4]^b2[6]^b2[7]^b2[8]^b2[11]^b2[12]^b2[13]^b2[14];//r0 + r4 + r6 + r7 + r8 + r11 + r12 + r13 + r14,       
         
         
         S13[15]=b7[2]^b7[4]^b7[6]^b7[7]^b7[8]^b7[9]^b7[10]^b7[11]^b7[13]^b7[14]^b7[15];           //   r2 + r4 + r6 + r7 + r8 + r9 + r10 + r11 + r13 + r14 + r15, 
         S13[14]=b7[4]^b7[6]^b7[8]^b7[10]^b7[11]^b7[15];//              r4 + r6 + r8 + r10 + r11 + r15,
         S13[13]=b7[1]^b7[2]^b7[3]^b7[5]^b7[6]^b7[7]^b7[8]^b7[10]^b7[11]^b7[12]^b7[13];//         r1 + r2 + r3 + r5 + r6 + r7 + r8 + r10 + r11 + r12 + r13,
         S13[12]=b7[2]^b7[4]^b7[7]^b7[9]^b7[10]^b7[11]^b7[14]^b7[15];//                    r2 + r4 + r7 + r9 + r10 + r11 + r14 + r15,
         S13[11]=b7[3]^b7[4]^b7[6]^b7[7]^b7[11]^b7[12]^b7[13]^b7[15];//             r3 + r4 + r6 + r7 + r11 + r12 + r13 + r15,
         S13[10]=b7[2]^b7[5]^b7[6]^b7[7]^b7[8]^b7[9]^b7[11]^b7[12]^b7[13]^b7[14]^b7[15];//     r2 + r5 + r6 + r7 + r8 + r9 + r11 + r12 + r13 + r14 + r15,
         S13[9]=b7[4]^b7[5]^b7[6]^b7[8]^b7[9]^b7[10]^b7[13]^b7[15];//         r4 + r5 + r6 + r8 + r9 + r10 + r13 + r15,
         S13[8]=b7[5]^b7[8]^b7[9];                                                          //          r5 + r8 + r9,
         S13[7]=b7[3]^b7[4]^b7[5]^b7[7]^b7[8]^b7[14];//                   r3 + r4 + r5 + r7 + r8 + r14,
         S13[6]=b7[3]^b7[4]^b7[8]^b7[10]^b7[11]^b7[12]^b7[15];//                  r3 + r4 + r8 + r10 + r11 + r12 + r15,
         S13[5]=b7[5]^b7[7]^b7[8]^b7[11]^b7[12]^b7[15];//                r5 + r7 + r8 + r11 + r12 + r15,
         S13[4]=b7[3]^b7[7]^b7[9]^b7[11]^b7[12]^b7[14]^b7[15];//          r3 + r7 + r9 + r11 + r12 + r14 + r15,
         S13[3]=b7[3]^b7[4]^b7[9]^b7[10]^b7[14]^b7[15];                     //              r3 + r4 + r9 + r10 + r14 + r15,
         S13[2]=b7[4]^b7[6]^b7[7]^b7[8]^b7[10]^b7[13]^b7[15];//               r4 + r6 + r7 + r8 + r10 + r13 + r15,
         S13[1]=b7[3]^b7[4]^b7[5]^b7[7]^b7[9]^b7[11]^b7[13]^b7[14];                                //   r3 + r4 + r5 + r7 + r9 + r11 + r13 + r14,
         S13[0]=b7[0]^b7[4]^b7[7]^b7[9]^b7[10]^b7[12]^b7[15];//     r0 + r4 + r7 + r9 + r10 + r12 + r15,    
         
         S14[15]=b4[2]^b4[4]^b4[5]^b4[6]^b4[8]^b4[13]^b4[14]^b4[15];//     r2 + r4 + r5 + r6 + r8 + r13 + r14 + r15,
         S14[14]=b4[1]^b4[2]^b4[3]^b4[5]^b4[7]^b4[8]^b4[10]^b4[11]^b4[12]^b4[15];//         r1 + r2 + r3 + r5 + r7 + r8 + r10 + r11 + r12 + r15,
         S14[13]=b4[4]^b4[5]^b4[8]^b4[14];//                             r4 + r5 + r8 + r14, 
         S14[12]=b4[2]^b4[5]^b4[7]^b4[8]^b4[9]^b4[10]^b4[12]^b4[13]^b4[14];//                       r2 + r5 + r7 + r8 + r9 + r10 + r12 + r13 + r14,
         S14[11]=b4[4]^b4[8]^b4[9]^b4[10]^b4[11]^b4[14]^b4[15];//                                       r4 + r8 + r9 + r10 + r11 + r14 + r15,
         S14[10]=b4[3]^b4[4]^b4[5]^b4[6]^b4[8]^b4[9]^b4[10]^b4[12]^b4[13]^b4[14]^b4[15];//         r3 + r4 + r5 + r6 + r8 + r9 + r10 + r12 + r13 + r14 + r15,
         S14[9]=b4[3]^b4[6]^b4[7]^b4[9]^b4[10]^b4[11]^b4[12];//                     r3 + r6 + r7 + r9 + r10 + r11 + r12, 
         S14[8]=b4[4]^b4[6]^b4[7]^b4[9]^b4[10]^b4[11]^b4[12];//                   r4 + r6 + r7 + r9 + r10 + r11 + r12,
         S14[7]=b4[3]^b4[5]^b4[7]^b4[8]^b4[10]^b4[13]^b4[14];//                   r3 + r5 + r7 + r8 + r10 + r13 + r14,
         S14[6]=b4[2]^b4[3]^b4[5]^b4[6]^b4[14]^b4[15];//                 r2 + r3 + r5 + r6 + r14 + r15,
         S14[5]=b4[3]^b4[5]^b4[6]^b4[8]^b4[9];//                     r3 + r5 + r6 + r8 + r9,
         S14[4]=b4[2]^b4[3]^b4[5]^b4[7]^b4[11]^b4[13]^b4[14]^b4[15];//                   r2 + r3 + r5 + r7 + r11 + r13 + r14 + r15,
         S14[3]=b4[2]^b4[3]^b4[6]^b4[13]^b4[15];                     //                                r2 + r3 + r6 + r13 + r15,    
         S14[2]=b4[3]^b4[5]^b4[6]^b4[7]^b4[9]^b4[10]^b4[11]^b4[14]^b4[15];//          r3 + r5 + r6 + r7 + r9 + r10 + r11 + r14 + r15,
         S14[1]=b4[2]^b4[6]^b4[7]^b4[8]^b4[9]^b4[11]^b4[12]^b4[13]^b4[14];              //                      r2 + r6 + r7 + r8 + r9 + r11 + r12 + r13 + r14,
         S14[0]=b4[0]^b4[3]^b4[6]^b4[8]^b4[10]^b4[11]^b4[13]^b4[14]^b4[15];//               r0 + r3 + r4 + r6 + r8 + r10 + r11 + r12 + r14 + r15,          
         
         S15[15]=b8[1]^b8[4]^b8[5]^b8[6]^b8[8]^b8[11]^b8[13]^b8[14]^b8[15];//     r1 + r4 + r5 + r6 + r7 + r8 + r11 + r12 + r13 + r14 + r15,
         S15[14]=b8[2]^b8[4]^b8[6]^b8[7]^b8[8]^b8[11]^b8[13]^b8[14];//                        r2 + r4 + r6 + r7 + r9 + r11 + r13 + r14,
         S15[13]=b8[3]^b8[8]^b8[10]^b8[11]^b8[12];//                                 r3 + r8 + r10 + r11 + r12,
         S15[12]=b8[3]^b8[4]^b8[5]^b8[6]^b8[8]^b8[10]^b8[13];//                        r3 + r4 + r5 + r6 + r8 + r10 + r13,
         S15[11]=b8[3]^b8[5]^b8[6]^b8[7]^b8[10]^b8[12]^b8[13]^b8[14];//                        r3 + r5 + r6 + r7 + r10 + r12 + r13 + r14,,
         S15[10]=b8[3]^b8[6]^b8[7]^b8[9]^b8[11]^b8[13]^b8[15];//                 r3 + r6 + r7 + r9 + r11 + r13 + r15,
         S15[9]=b8[2]^b8[3]^b8[4]^b8[5]^b8[7]^b8[12]^b8[15];//                          r2 + r3 + r4 + r5 + r7 + r12 + r15,
         S15[8]=b8[3]^b8[5]^b8[7]^b8[9]^b8[10]^b8[11]^b8[15];//                      r3 + r5 + r7 + r9 + r10 + r11 + r15,
         S15[7]=b8[5]^b8[6]^b8[7]^b8[8]^b8[8]^b8[9]^b8[11]^b8[13]^b8[14];//                      r5 + r6 + r7 + r8 + r9 + r11 + r13 + r14,
         S15[6]=b8[3]^b8[4]^b8[7]^b8[8]^b8[9]^b8[10]^b8[11]^b8[12]^b8[13]^b8[15];//                  r3 + r4 + r7 + r8 + r9 + r10 + r11 + r12 + r13 + r15,
         S15[5]=b8[2]^b8[3]^b8[5]^b8[9]^b8[10]^b8[11]^b8[12]^b8[13]^b8[14];//                       r2 + r3 + r5 + r9 + r10 + r11 + r12 + r13 + r14, 
         S15[4]=b8[2]^b8[6]^b8[8]^b8[11]^b8[13]^b8[14];//                        r2 + r6 + r8 + r11 + r13 + r14, 
         S15[3]=b8[2]^b8[5]^b8[6]^b8[7]^b8[8]^b8[9]^b8[10]^b8[13]^b8[14]; //                    r2 + r5 + r6 + r7 + r8 + r9 + r10 + r13 + r14, 
         S15[2]=b8[3]^b8[5]^b8[6]^b8[7]^b8[9]^b8[10]^b8[11]^b8[14]^b8[15];//          r3 + r5 + r6 + r7 + r9 + r10 + r11 + r14 + r15,
         S15[1]=b8[2]^b8[3]^b8[4]^b8[5]^b8[9]^b8[10];   //              r2 + r3 + r4 + r5 + r9 + r10,
         S15[0]=b8[0]^b8[2]^b8[6]^b8[7]^b8[13]^b8[14];//                r0 + r2 + r6 + r7 + r13 + r14,        
         
         S16[15]=b1[3]^b1[5]^b1[6]^b1[7]^b1[9]^b1[10]^b1[15];//r3 + r5 + r6 + r7 + r9 + r10 + r15,
         S16[14]=b1[7]^b1[8]^b1[9]^b1[10]^b1[13]^b1[14]^b1[15];//               r7 + r8 + r9 + r10 + r13 + r14 + r15,
         S16[13]=b1[3]^b1[5]^b1[7]^b1[8]^b1[9]^b1[12]^b1[13];//            r3 + r5 + r7 + r8 + r9 + r12 + r13,
         S16[12]=b1[3]^b1[4]^b1[5]^b1[6]^b1[7]^b1[8]^b1[9]^b1[12]^b1[13];//       r3 + r4 + r5 + r6 + r7 + r8 + r9 + r12 + r13,
         S16[11]=b1[3]^b1[5]^b1[7]^b1[8]^b1[9]^b1[11]^b1[12];//          r3 + r5 + r7 + r8 + r9 + r11 + r12,
         S16[10]=b1[2]^b1[3]^b1[6]^b1[7]^b1[8]^b1[10]^b1[14]^b1[15];//     r2 + r3 + r6 + r7 + r8 + r10 + r14 + r15, 
         S16[9]=b1[4]^b1[10]^b1[11]^b1[12]^b1[13]^b1[15];//                         r4 + r10 + r11 + r12 + r13 + r15,
         S16[8]=b1[3]^b1[4]^b1[10]^b1[12]^b1[13]^b1[14]^b1[15];//    r3 + r4 + r10 + r12 + r13 + r14 + r15,
         S16[7]=b1[3]^b1[4]^b1[6]^b1[7]^b1[8]^b1[9]^b1[12]^b1[14];//        r3 + r4 + r6 + r7 + r8 + r9 + r12 + r14,
         S16[6]=b1[2]^b1[4]^b1[5]^b1[6]^b1[9]^b1[10]^b1[11]^b1[12]^b1[14];//  r2 + r4 + r5 + r6 + r9 + r10 + r11 + r12 + r14,
         S16[5]=b1[1]^b1[3]^b1[5]^b1[6]^b1[7];//          r1 + r3 + r5 + r6 + r7,
         S16[4]=b1[2]^b1[3]^b1[4]^b1[6]^b1[8]^b1[11]^b1[13]^b1[14];//               r2 + r3 + r4 + r6 + r8 + r11 + r13 + r14,,
         S16[3]=b1[1]^b1[3]^b1[8]^b1[9]^b1[10]^b1[12]^b1[13]^b1[15];// r1 + r3 + r8 + r9 + r10 + r12 + r13 + r15,
         S16[2]=b1[1]^b1[3]^b1[5]^b1[13]^b1[15];//          r1 + r3 + r5 + r13 + r15,
         S16[1]=b1[5]^b1[6]^b1[7]^b1[10]^b1[11]^b1[12]^b1[15]; //                     r5 + r6 + r7 + r10 + r11 + r12 + r15,
         S16[0]=b1[0]^b1[1]^b1[2]^b1[3]^b1[4]^b1[5]^b1[6]^b1[7]^b1[9]^b1[11]^b1[15];// r0 + r1 + r2 + r3 + r4 + r5 + r6 + r7 + r9 + r11 + r15,
        
         S17[15]=b9[3]^b9[8]^b9[9]^b9[11]^b9[12]^b9[14];// r3 + r8 + r9 + r11 + r12 + r14,
         S17[14]=b9[3]^b9[7]^b9[10]^b9[12]^b9[14];//               r3 + r7 + r10 + r12 + r14,
         S17[13]=b9[3]^b9[4]^b9[6]^b9[9]^b9[14];//                 r3 + r4 + r6 + r9 + r14,
         S17[12]=b9[2]^b9[4]^b9[6]^b9[7]^b9[8]^b9[10]^b9[11]^b9[14];//      r2 + r4 + r6 + r7 + r8 + r10 + r11 + r14,
         S17[11]=b9[3]^b9[4]^b9[5]^b9[6]^b9[7]^b9[10]^b9[13];//          r3 + r4 + r5 + r6 + r7 + r10 + r13,
         S17[10]=b9[3]^b9[4]^b9[5]^b9[7]^b9[8]^b9[10]^b9[12];//      r3 + r4 + r5 + r7 + r8 + r9 + r10 + r12, 
         S17[9]=b9[5]^b9[12];//                         r5 + r12,
         S17[8]=b9[2]^b9[3]^b9[4]^b9[6]^b9[8]^b9[9]^b9[11]^b9[12]^b9[14];//    r2 + r3 + r4 + r6 + r8 + r9 + r11 + r12 + r14,
         S17[7]=b9[5]^b9[6]^b9[8]^b9[9]^b9[11]^b9[13]^b9[14]^b9[15];//         r5 + r6 + r8 + r9 + r11 + r13 + r14 + r15,
         S17[6]=b9[1]^b9[2]^b9[3]^b9[5]^b9[6]^b9[8]^b9[11]^b9[14]^b9[15];//  r1 + r2 + r3 + r5 + r6 + r8 + r11 + r14 + r15,
         S17[5]=b9[3]^b9[4]^b9[5]^b9[6]^b9[7]^b9[8]^b9[10]^b9[12]^b9[13];//         r3 + r4 + r5 + r6 + r7 + r8 + r10 + r12 + r13,
         S17[4]=b9[1]^b9[3]^b9[4]^b9[5]^b9[6]^b9[7]^b9[9]^b9[13]^b9[14];//            r1 + r3 + r4 + r5 + r6 + r7 + r9 + r13 + r14,
         S17[3]=b9[1]^b9[4]^b9[6]^b9[8]^b9[9]^b9[11]^b9[12]^b9[13]^b9[14];// r1 + r4 + r6 + r8 + r9 + r11 + r12 + r13 + r14,
         S17[2]=b9[2]^b9[4]^b9[7]^b9[8]^b9[9]^b9[12]^b9[14]^b9[15];//              r2 + r4 + r7 + r8 + r9 + r12 + r14 + r15,
         S17[1]=b9[1]^b9[5]^b9[7]^b9[11]^b9[13]^b9[14]; //                  r1 + r5 + r7 + r11 + r13 + r14,
         S17[0]=b9[0]^b9[3]^b9[4]^b9[5]^b9[6]^b9[9]^b9[10]^b9[15];//  r0 + r3 + r4 + r5 + r6 + r9 + r10 + r15,
         
          S18[15]=b5[4]^b5[5]^b5[8]^b5[10]^b5[11]^b5[15];                         //      r4 + r5 + r8 + r10 + r11 + r15,
          S18[14]=b5[2]^b5[3]^b5[4]^b5[5]^b5[6]^b5[8]^b5[11]^b5[13];//              r2 + r3 + r4 + r5 + r6 + r8 + r11 + r13,
          S18[13]=b5[3]^b5[6]^b5[8]^b5[10]^b5[11]^b5[13]^b5[14];//         r3 + r6 + r8 + r10 + r11 + r13 + r14,
          S18[12]=b5[4]^b5[5]^b5[6]^b5[7]^b5[8]^b5[9]^b5[11]^b5[12];//        r4 + r5 + r6 + r7 + r8 + r9 + r11 + r12,
          S18[11]=b5[3]^b5[5]^b5[6]^b5[7]^b5[8]^b5[9]^b5[13]^b5[15];//               r3 + r5 + r6 + r7 + r8 + r9 + r13 + r15,
          S18[10]=b5[2]^b5[5]^b5[6]^b5[7]^b5[9]^b5[10]^b5[13]^b5[15];//                 r2 + r5 + r6 + r7 + r9 + r10 + r13 + r15,
          S18[9]=b5[3]^b5[4]^b5[5]^b5[6]^b5[7]^b5[11]^b5[13]^b5[15];//              r3 + r4 + r5 + r6 + r7 + r11 + r13 + r15,
          S18[8]=b5[2]^b5[3]^b5[4]^b5[6]^b5[7]^b5[9]^b5[10]^b5[11]^b5[13];//          r2 + r3 + r4 + r6 + r7 + r9 + r10 + r11 + r13,
          S18[7]=b5[1]^b5[4]^b5[6]^b5[8]^b5[15];//                      r1 + r4 + r6 + r8 + r15,
          S18[6]=b5[3]^b5[5]^b5[6]^b5[8]^b5[9]^b5[12];//                      r3 + r5 + r6 + r8 + r9 + r12,
          S18[5]=b5[1]^b5[4]^b5[7]^b5[10]^b5[15];//              r1 + r4 + r7 + r10 + r15,
          S18[4]=b5[1]^b5[2]^b5[9]^b5[10]^b5[13]^b5[14]^b5[15];//                   r1 + r2 + r9 + r10 + r13 + r14 + r15,
          S18[3]=b5[3]^b5[5]^b5[8]^b5[9]^b5[14]^b5[15];//                   r3 + r5 + r8 + r9 + r14 + r15,
          S18[2]=b5[1]^b5[4]^b5[5]^b5[6]^b5[7]^b5[9]^b5[11]^b5[12]^b5[14];//      r1 + r4 + r5 + r6 + r7 + r9 + r11 + r12 + r14,
          S18[1]=b5[3]^b5[4]^b5[6]^b5[9]^b5[11]^b5[12]^b5[13]^b5[15]; //              r3 + r4 + r6 + r7 + r9 + r11 + r12 + r13 + r15,
          S18[0]=b5[0]^b5[3]^b5[4]^b5[5]^b5[8]^b5[9]^b5[12]^b5[13]^b5[14];//             r0 + r3 + r4 + r5 + r8 + r9 + r12 + r13 + r14,
         
         
         S19[15]=b10[5]^b10[6]^b10[7]^b10[8]^b10[9]^b10[11]^b10[13]^b10[15];                         //r5 + r6 + r7 + r8 + r9 + r10 + r11 + r13 + r15,
         S19[14]=b10[3]^b10[5]^b10[6]^b10[8]^b10[11]^b10[12];//                 r3 + r5 + r6 + r8 + r11 + r12,
         S19[13]=b10[4]^b10[6]^b10[9]^b10[11]^b10[14];//                r4 + r6 + r9 + r11 + r14,
         S19[12]=b10[2]^b10[3]^b10[4]^b10[6]^b10[7]^b10[8]^b10[9]^b10[12];//            r2 + r3 + r4 + r6 + r7 + r8 + r9 + r12,
         S19[11]=b10[3]^b10[4]^b10[5]^b10[9]^b10[10]^b10[12]^b10[13]^b10[14]^b10[15];//               r3 + r4 + r5 + r9 + r10 + r12 + r13 + r14 + r15,
         S19[10]=b10[2]^b10[10]^b10[11]^b10[12];//                         r2 + r10 + r11 + r12,
         S19[9]=b10[3]^b10[4]^b10[5]^b10[6]^b10[7]^b10[8]^b10[10]^b10[11]^b10[15];//          r3 + r4 + r5 + r6 + r7 + r8 + r10 + r11 + r15,
         S19[8]=b10[1]^b10[4]^b10[12]^b10[13];//                 r1 + r4 + r12 + r13,
         S19[7]=b10[4]^b10[6]^b10[7]^b10[8]^b10[10]^b10[12]^b10[14];//                           r4 + r6 + r7 + r8 + r10 + r12 + r14,
         S19[6]=b10[1]^b10[2]^b10[5]^b10[6]^b10[8]^b10[9]^b10[10]^b10[14]^b10[15];//                       r1 + r2 + r5 + r6 + r8 + r9 + r10 + r14 + r15,
         S19[5]=b10[1]^b10[2]^b10[3]^b10[5]^b10[6]^b10[7]^b10[10]^b10[11]^b10[12]^b10[14]^b10[15];//               r1 + r2 + r3 + r5 + r6 + r7 + r10 + r11 + r12 + r14 + r15,
         S19[4]=b10[6]^b10[8]^b10[11]^b10[12]^b10[13]^b10[15];//                           r6 + r8 + r11 + r12 + r13 + r15,
         S19[3]=b10[1]^b10[2]^b10[3]^b10[5]^b10[6]^b10[7]^b10[8]^b10[11]^b10[14]^b10[15];//                  r1 + r2 + r3 + r5 + r6 + r7 + r8 + r11 + r14 + r15,
         S19[2]=b10[2]^b10[3]^b10[5]^b10[10]^b10[12]^b10[13]^b10[14]^b10[15];//        r2 + r3 + r5 + r10 + r12 + r13 + r14 + r15,
         S19[1]=b10[3]^b10[5]^b10[6]^b10[7]^b10[9]^b10[13]^b10[14]^b10[15]; //             r3 + r5 + r6 + r7 + r9 + r13 + r14 + r15,
         S19[0]=b10[0]^b10[2]^b10[3]^b10[4]^b10[5]^b10[6]^b10[7]^b10[13];//            r0 + r2 + r3 + r4 + r5 + r6 + r7 + r13,
         
         
         S20[15]=b3[3]^b3[4]^b3[6]^b3[8]^b3[9]^b3[10]^b3[12]^b3[14]^b3[15];//                 r3 + r4 + r6 + r8 + r9 + r10 + r12 + r14 + r15,
         S20[14]=b3[2]^b3[3]^b3[5]^b3[7]^b3[8]^b3[10]^b3[12]^b3[15];//         r2 + r3 + r5 + r7 + r8 + r10 + r12 + r15,
         S20[13]=b3[4]^b3[6]^b3[9]^b3[14];//       r4 + r6 + r9 + r14,
         S20[12]=b3[2]^b3[3]^b3[4]^b3[6]^b3[7]^b3[13]^b3[14]^b3[15];//      r2 + r3 + r4 + r6 + r7 + r13 + r14 + r15,
         S20[11]=b3[4]^b3[5]^b3[6]^b3[7]^b3[10]^b3[13]^b3[15];                    //                   r4 + r5 + r6 + r7 + r10 + r13 + r15,
         S20[10]=b3[5]^b3[7]^b3[8]^b3[9]^b3[10]^b3[11]^b3[12]^b3[14]^b3[15];//             r5 + r7 + r8 + r9 + r10 + r11 + r12 + r14 + r15,
         S20[9]=b3[1]^b3[5]^b3[7]^b3[8]^b3[12]^b3[15];//                         r1 + r5 + r7 + r8 + r12 + r15,
         S20[8]=b3[2]^b3[3]^b3[7]^b3[8]^b3[9]^b3[12];//                                       r2 + r3 + r7 + r8 + r9 + r12,
         S20[7]=b3[1]^b3[2]^b3[7]^b3[13]^b3[15];//                        r1 + r2 + r7 + r13 + r15,
         S20[6]=b3[1]^b3[4]^b3[5]^b5[6]^b3[8]^b3[10]^b3[11]^b3[14]^b3[15];//                r1 + r4 + r5 + r6 + r8 + r10 + r11 + r14 + r15,
         S20[5]=b3[2]^b3[3]^b3[4]^b3[5]^b3[6]^b3[9]^b3[10]^b3[13];//              r2 + r3 + r4 + r5 + r6 + r9 + r10 + r13,
         S20[4]=b3[1]^b3[2]^b3[5]^b3[9]^b3[11];//                                r1 + r2 + r5 + r9 + r11,
         S20[3]=b3[6]^b3[8]^b3[10]^b3[11]^b3[12];//                      r6 + r8 + r10 + r11 + r12,
         S20[2]=b3[2]^b3[4]^b3[5]^b3[6]^b3[7]^b3[10]^b3[11]^b3[12]^b3[15];//  r2 + r4 + r5 + r6 + r7 + r10 + r11 + r12 + r15, 
         S20[1]=b3[3]^b3[4]^b3[8]^b3[10]^b3[12]^b3[14]; //                    r3 + r4 + r8 + r10 + r12 + r14,
         S20[0]=b3[0]^b3[4]^b3[5]^b3[7]^b3[10]^b3[11]^b3[12];//                   r0 + r4 + r5 + r7 + r10 + r11 + r12,  
         
         S21[15]=b11[3]^b11[4]^b11[7]^b11[10]^b11[11]^b11[14];//               r3 + r4 + r5 + r7 + r10 + r11 + r14,
         S21[14]=b11[2]^b11[5]^b11[7]^b11[8]^b11[9]^b11[10]^b11[11]^b11[13]^b11[14]^b11[15];//            r2 + r5 + r7 + r8 + r9 + r10 + r11 + r13 + r14 + r15,
         S21[13]=b11[11]^b11[12]^b11[13];//            r11 + r12 + r13,
         S21[12]=b11[6]^b11[8]^b11[13]^b11[14];//              r6 + r8 + r13 + r14,
         S21[11]=b11[3]^b11[5]^b11[6]^b11[10]^b11[11];                    //                   r3 + r5 + r6 + r10 + r11,
         S21[10]=b11[1]^b11[2]^b11[4]^b11[5]^b11[6]^b11[7]^b11[8]^b11[9]^b11[10]^b11[11]^b11[13]^b11[15];//         r1 + r2 + r4 + r5 + r6 + r7 + r8 + r9 + r10 + r11 + r13 + r15,
         S21[9]=b11[2]^b11[4]^b11[5]^b11[6]^b11[7]^b11[8]^b11[9]^b11[14];//                           r2 + r4 + r5 + r6 + r7 + r8 + r9 + r14,
         S21[8]=b11[1]^b11[3]^b11[4]^b11[5]^b11[6]^b11[8]^b11[9]^b11[11]^b11[13]^b11[14];//                             r1 + r3 + r4 + r5 + r6 + r8 + r9 + r11 + r13 + r14,
         S21[7]=b11[1]^b11[2]^b11[3]^b11[5]^b11[7]^b11[11];//                              r1 + r2 + r3 + r5 + r7 + r11,
         S21[6]=b11[2]^b11[3]^b11[4]^b11[5]^b11[9]^b11[11]^b11[13]^b11[14];//          r2 + r3 + r4 + r5 + r9 + r10 + r11 + r13 + r14,
         S21[5]=b11[1]^b11[2]^b11[3]^b11[4]^b11[5]^b11[6]^b11[9]^b11[11]^b11[13]^b11[14];//             r1 + r2 + r3 + r4 + r5 + r6 + r9 + r11 + r13 + r14,
         S21[4]=b11[2]^b11[3]^b11[9]^b11[10]^b11[11]^b11[12]^b11[15];//                                   r2 + r3 + r9 + r10 + r11 + r12 + r15,
         S21[3]=b11[2]^b11[3]^b11[4]^b11[7]^b11[10]^b11[11]^b11[12];//                         r2 + r3 + r4 + r7 + r10 + r11 + r12,
         S21[2]=b11[2]^b11[3]^b11[4]^b11[5]^b11[6]^b11[10]^b11[12]^b11[13]^b11[14];//    r2 + r3 + r4 + r5 + r6 + r10 + r12 + r13 + r14,
         S21[1]=b11[3]^b11[4]^b11[6]^b11[7]^b11[8]^b11[9]^b11[11]; //                          r3 + r4 + r6 + r7 + r8 + r9 + r11,
         S21[0]=b11[0]^b11[2]^b11[4]^b11[5]^b11[7]^b11[8]^b11[10]^b11[12]^b11[15];//                    r0 + r2 + r4 + r5 + r7 + r8 + r10 + r12 + r15,
         
         S22[15]=b6[5]^b6[6]^b6[9]^b6[12]^b6[14];//             r5 + r6 + r9 + r12 + r14,
         S22[14]=b6[3]^b6[4]^b6[5]^b6[6]^b6[7]^b6[9]^b6[14]^b6[15];//            r3 + r4 + r5 + r6 + r7 + r9 + r14 + r15,
         S22[13]=b6[4]^b6[5]^b6[9]^b6[15];//                     r4 + r5 + r9 + r15,
         S22[12]=b6[1]^b6[2]^b6[3]^b6[4]^b6[6]^b6[10]^b6[12]^b6[13]^b6[14]^b6[15];//                    r2 + r4 + r5 + r9 + r11 + r13 + r14 + r15,
         S22[11]=b6[1]^b6[2]^b6[3]^b6[5]^b6[6]^b6[7]^b6[8]^b6[11]^b6[12]^b6[14]^b6[15];                    //               r1 + r2 + r3 + r5 + r6 + r7 + r8 + r11 + r12 + r14 + r15,
         S22[10]=b6[3]^b6[4]^b6[5]^b6[10]^b6[11]^b6[13];//              r3 + r4 + r5 + r10 + r11 + r13,
         S22[9]=b6[1]^b6[2]^b6[3]^b6[4]^b6[5]^b6[7]^b6[8]^b6[9]^b6[12]^b6[14]^b6[15];//                      r1 + r2 + r3 + r4 + r5 + r7 + r8 + r9 + r12 + r14 + r15,
         S22[8]=b6[1]^b6[2]^b6[3]^b6[4]^b6[5]^b6[6]^b6[7]^b6[9]^b6[15];//                      r1 + r2 + r3 + r4 + r5 + r6 + r7 + r9 + r15,
         S22[7]=b6[2]^b6[4]^b6[13]^b6[14]^b6[15];//                                  r2 + r4 + r13 + r14 + r15,
         S22[6]=b6[1]^b6[2]^b6[3]^b6[6]^b6[8]^b6[10]^b6[11]^b6[13]^b6[15];//             r1 + r2 + r3 + r6 + r8 + r10 + r11 + r13 + r15,
         S22[5]=b6[5]^b6[12]^b6[15];//                  r5 + r12 + r15,
         S22[4]=b6[2]^b6[4]^b6[5]^b6[7]^b6[8]^b6[10]^b6[13]^b6[14]^b6[15];//                              r2 + r4 + r5 + r7 + r8 + r10 + r13 + r14 + r15,
         S22[3]=b6[2]^b6[4]^b6[10]^b6[11]^b6[12];//                          r2 + r4 + r10 + r11 + r12,
         S22[2]=b6[3]^b6[5]^b6[7]^b6[9]^b6[10]^b6[12]^b6[14];//          r3 + r5 + r7 + r9 + r10 + r12 + r14,
         S22[1]=b6[6]^b6[7]^b6[8]^b6[9]^b6[11]^b6[14]; //                            r6 + r7 + r8 + r9 + r11 + r14,
         S22[0]=b6[0]^b6[2]^b6[5]^b6[6]^b6[7]^b6[8]^b6[10]^b6[11]^b6[12]^b6[13]^b6[15];//              r0 + r2 + r5 + r6 + r7 + r8 + r10 + r11 + r12 + r13 + r15,
         
         
         S23[15]=b12[5]^b12[7]^b12[12];//                 r5 + r7 + r12]
         S23[14]=b12[2]^b12[3]^b12[4]^b12[5]^b12[6]^b12[8]^b12[10]^b12[11]^b12[13];//           r2 + r3 + r4 + r5 + r6 + r8 + r10 + r11 + r13]
         S23[13]=b12[2]^b12[3]^b12[4]^b12[5]^b12[9]^b12[10]^b12[15];//                        r2 + r3 + r4 + r5 + r9 + r10 + r12 + r13]
         S23[12]=b12[1]^b12[3]^b12[4]^b12[6]^b12[8]^b12[9]^b12[10]^b12[15];//                       r1 + r3 + r4 + r6 + r8 + r9 + r10 + r15]
         S23[11]=b12[2]^b12[3]^b12[4]^b12[7]^b12[9]^b12[12]^b12[13]^b12[14]^b12[15];                    //              r2 + r3 + r4 + r7 + r9 + r12 + r13 + r14 + r15]
         S23[10]=b12[1]^b12[2]^b12[5]^b12[6]^b12[7]^b12[10]^b12[13]^b12[14];//                  r1 + r2 + r5 + r6 + r7 + r10 + r13 + r14]
         S23[9]=b12[1]^b12[2]^b12[3]^b12[6]^b12[7]^b12[8]^b12[12]^b12[13]^b12[15];//                    r1 + r2 + r3 + r6 + r7 + r8 + r10 + r12 + r13 + r15]
         S23[8]=b12[2]^b12[4]^b12[5]^b12[6]^b12[9]^b12[12]^b12[13]^b12[14];//                      r2 + r4 + r5 + r6 + r9 + r12 + r13 + r14]
         S23[7]=b12[1]^b12[5]^b12[6]^b12[7]^b12[9]^b12[10];//                                         r1 + r5 + r6 + r7 + r9 + r10]
         S23[6]=b12[2]^b12[3]^b12[4]^b12[5]^b12[6]^b12[10]^b12[12]^b12[13]^b12[14];//                r2 + r3 + r4 + r5 + r6 + r10 + r12 + r13 + r14]
         S23[5]=b12[2]^b12[3]^b12[6]^b12[7]^b12[8]^b12[10]^b12[11]^b12[13]^b12[14]^b12[15];//                  r2 + r3 + r6 + r7 + r8 + r10 + r11 + r13 + r14 + r15]
         S23[4]=b12[3]^b12[5]^b12[7]^b12[8]^b12[10]^b12[11]^b12[12]^b12[14]^b12[15];//                           r3 + r5 + r7 + r8 + r10 + r11 + r12 + r14 + r15]
         S23[3]=b12[3]^b12[5]^b12[6]^b12[7]^b12[9]^b12[10]^b12[11]^b12[14];//                         r3 + r5 + r6 + r7 + r9 + r10 + r11 + r14]
         S23[2]=b12[2]^b12[9]^b12[10]^b12[12]^b12[15];//              r2 + r9 + r10 + r12 + r15]
         S23[1]=b12[3]^b12[4]^b12[5]^b12[6]^b12[8]^b12[9]^b12[11]^b12[12]^b12[13]^b12[14]^b12[15]; //          r3 + r4 + r5 + r6 + r8 + r9 + r11 + r12 + r13 + r14 + r15]
         S23[0]=b12[0]^b12[4]^b12[5]^b12[7]^b12[10]^b12[12];//                r0 + r4 + r5 + r7 + r10 + r12]
        
        
                  
                  
         
         
         
         
         
         
         
         
         
         
  /*       S[1]=S1;    
         S[2]=S2;   
         S[3]=S3;   
         S[4]=S4;   
         S[5]=S5;   
         S[6]=S6;   
         S[7]=S7;   
         S[8]=S8;   
         S[9]=S9;   
         S[10]=S10;   
         S[11]=S11;   
         S[12]=S12;   
         S[13]=S13;   
         S[14]=S14;   
         S[15]=S15;   
         S[16]=S16;   
         S[17]=S17;   
         S[18]=S18;   
         S[19]=S19;   
         S[20]=S20;   
         S[21]=S21;   
         S[22]=S22;   
         S[23]=S23;   */
         
              
                  
                  
                  
                  end
                  
          /*     if(count>16200)
                begin
                count=16208;            //2019.05.26  �ɸ�ֵΪ��ĳ�16208
         
                
                enableBM=1;
                     
                i=0;
                j=191;
                end     */
              end
          
    /*              always@(posedge CLK)
              begin
              if (count<=16008)
                    Cfront[count-1]<=R;
              end    
      */
      always@(posedge CLK)
      if((count>16200)&&(count<=16201))
                      begin
                      count=count+1;            //2019.05.26  �ɸ�ֵΪ��ĳ�16208
                            
                     enableBM=1;
                           
                      i=0;
                      j=191;
                      end 
        
        always@(posedge CLK)
                            if(count==16202)
                                            begin
                                            count=count+1;            //2019.05.26  �ɸ�ֵΪ��ĳ�16208
                                                  
                                           enableBM=1;
                                                 
                                            i=0;
                                            j=191;
                                            end 
                      

endmodule
